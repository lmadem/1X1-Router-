// Code your testbench here
// or browse Examples
`include "top.sv"
`include "router_if.sv"
`include "program_router_tb.sv"
