//test_sa2 : This test is to send the stimulus from a single source port to various destination ports (SA2 -> DA*)

class test_sa2 extends uvm_test;
  //Register test_sa2 into factory
  `uvm_component_utils(test_sa2);
  
  //Instantiate environment component
  environment env;
  
  //virtual interface
  virtual router_if vif;
  
  //custom constructor
  function new (string name = "test_sa2", uvm_component parent);
    super.new(name, parent);
  endfunction
  
  //extern methods
  extern virtual function void build_phase(uvm_phase phase);
  extern virtual function void start_of_simulation_phase(uvm_phase phase);
  extern virtual task main_phase(uvm_phase phase);

endclass	

//build_phase to construct child components
function void test_sa2::build_phase(uvm_phase phase);
  super.build_phase(phase);
  
  //Construct object for environment
  env = environment::type_id::create("env", this);
  
  //Below shown all are environment(testbench) configurations
  //Get the physical interface from program block
  uvm_config_db#(virtual router_if)::get(this, "", "vif", vif);
  
  //set the test name for readability in the environment
  uvm_config_db#(string)::set(this, "env.*", "test_name", get_type_name());
  
  //below are to set the physical interface to child components (drvr,iMon and oMon) 
  //Set the physical interface to Driver
  uvm_config_db#(virtual router_if.tb_mod_port)::set(this, "env.m_agent", "drvr_if", vif.tb_mod_port);
  
  //Set the physical interface to Input Monitor
  uvm_config_db#(virtual router_if.tb_mon)::set(this, "env.m_agent", "iMon_if", vif.tb_mon);
  
  //Set the physical interface to Output Monitor
  uvm_config_db#(virtual router_if.tb_mon)::set(this, "env.s_agent", "oMon_if", vif.tb_mon);
  
  //Set the number of packets to be generated by sequence
  uvm_config_db#(int)::set(this, "env.*", "item_count", 10);
  
  //Below shown settings are to configure sequencer to execute particular sequence in a particular phase
  
  //configure sequencer to execute reset_sequence in reset_phase of sequencer
  uvm_config_db#(uvm_object_wrapper)::set(this, "env.m_agent.seqr.reset_phase", "default_sequence", reset_sequence::get_type());
  
  //configure sequencer to execute config_sequence in configure_phase of sequencer
  uvm_config_db#(uvm_object_wrapper)::set(this, "env.m_agent.seqr.configure_phase", "default_sequence", config_sequence::get_type());
  
  //configure sequencer to execute sa2_sequence in main_phase of sequencer
  uvm_config_db#(uvm_object_wrapper)::set(this, "env.m_agent.seqr.main_phase", "default_sequence", sa2_sequence::get_type());
  
  
  //configure sequencer to execute shutdown_sequence in shutdown_phase of sequencer
  uvm_config_db#(uvm_object_wrapper)::set(this, "env.m_agent.seqr.shutdown_phase", "default_sequence", shutdown_sequence::get_type());

endfunction

//start_of_simulation_phase to print testbench topology
function void test_sa2::start_of_simulation_phase(uvm_phase phase);
  super.start_of_simulation_phase(phase);
  //Print testbench topology
  uvm_root::get().print_topology();
  
  //Print factory override information
  uvm_factory::get().print();

endfunction

//main_phase to set drain_time
task test_sa2::main_phase(uvm_phase phase);
  uvm_objection objection;
  super.main_phase(phase);
  
  //Get the phase objection object
  objection = phase.get_objection();
  
  //Set the Drain time..
  objection.set_drain_time(this, 25000ns);
  
  //The drain time is the amount of time to wait once all objections have been dropped
  
endtask



